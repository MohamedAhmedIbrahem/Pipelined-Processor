
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FETCH_DC_BUFFER IS
    PORT(
        CLK, RST, IR_HIGH_EN, IR_LOW_EN : IN  STD_LOGIC;
        P_TAKEN_IN      		: IN  STD_LOGIC;
	P_TAKEN_OUT 			: OUT STD_LOGIC;
        PC_KEY_IN          		: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        PC_KEY_OUT            		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        IR_FETCH             		: IN  STD_LOGIC_VECTOR(0 TO 15);
        IR_HIGH_OUT            		: OUT STD_LOGIC_VECTOR(0 TO 15);
        IR_LOW_OUT           		: OUT STD_LOGIC_VECTOR(0 TO 15)
    );
END ENTITY;

ARCHITECTURE arch OF FETCH_DC_BUFFER IS
	COMPONENT IR_HIGH IS
    	PORT(
        	CLK, RST, EN    : IN  STD_LOGIC;
        	Din             : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
       		Dout            : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    	);
	END COMPONENT;

	COMPONENT IR_LOW IS
    	PORT(
        	CLK, RST, EN    : IN  STD_LOGIC;
        	Din             : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
        	Dout            : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    	);
	END COMPONENT;
	COMPONENT PREDICTION_REG IS
    	PORT(
        	CLK, RST, EN    	: IN  STD_LOGIC;
        	P_TAKEN_IN      	: IN  STD_LOGIC;
		P_TAKEN_OUT 		: OUT STD_LOGIC;
        	PC_KEY_IN          	: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        	PC_KEY_OUT            	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    	);
	END COMPONENT;
	SIGNAL IR_High_Reg, IR_Low_Reg : STD_LOGIC_VECTOR(0 TO 15);
BEGIN
    	IR_High_Reg <= IR_FETCH WHEN IR_FETCH(0) = '0' ELSE (OTHERS => '0');
    	IR_Low_Reg <= IR_FETCH WHEN IR_FETCH(0) = '1' ELSE (OTHERS => '0');

	IR_REG_HIGH : IR_HIGH PORT MAP (CLK, RST, IR_HIGH_EN, IR_High_Reg, IR_HIGH_OUT);
	IR_REG_LOW : IR_LOW PORT MAP (CLK, RST, IR_LOW_EN, IR_Low_Reg, IR_LOW_OUT);
	PREDICT_REG : PREDICTION_REG PORT MAP (CLK, RST, IR_HIGH_EN, P_TAKEN_IN, P_TAKEN_OUT, PC_KEY_IN, PC_KEY_OUT);

END ARCHITECTURE;