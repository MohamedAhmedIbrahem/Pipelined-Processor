LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PREDICTION_REG IS
    PORT(
        CLK, RST, EN    	: IN  STD_LOGIC;
        P_TAKEN_IN      	: IN  STD_LOGIC;
	P_TAKEN_OUT 		: OUT STD_LOGIC;
        PC_KEY_IN          	: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        PC_KEY_OUT            	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch OF PREDICTION_REG IS
COMPONENT RISING_EDGE_REG IS
    GENERIC(Size: INTEGER := 32);
    PORT(
        CLK, RST, EN    : IN  STD_LOGIC;
        Din             : IN  STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
        Dout            : OUT STD_LOGIC_VECTOR(Size-1 DOWNTO 0)
    );
END COMPONENT;
BEGIN
    REG : RISING_EDGE_REG GENERIC MAP (4) PORT MAP (CLK => CLK , RST => RST , EN => EN , Din => PC_KEY_IN , Dout => PC_KEY_OUT);
	PROCESS(CLK, RST)
    BEGIN
        IF RISING_EDGE(CLK) THEN 
            IF RST='1' THEN
                P_TAKEN_OUT <= '0';
            ELSIF EN='1' THEN
                P_TAKEN_OUT <= P_TAKEN_IN;
            END IF;
        END IF;
    END PROCESS;
END ARCHITECTURE;