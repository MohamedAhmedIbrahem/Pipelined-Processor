LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PREDICTION_REG IS
    GENERIC(Size: INTEGER := 5);
    PORT(
        CLK, RST, EN    : IN  STD_LOGIC;
        P_TAKEN         : IN  STD_LOGIC;
        PC_KEY          : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Dout            : OUT STD_LOGIC_VECTOR(Size-1 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch OF PREDICTION_REG IS
SIGNAL Din : STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
BEGIN
    Din <= PC_KEY & P_TAKEN;
    REG : ENTITY work.RISING_EDGE_REG GENERIC MAP (Size) PORT MAP (CLK => CLK , RST => RST , EN => EN , Din => Din , Dout => Dout);
END ARCHITECTURE;